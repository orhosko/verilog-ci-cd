module our;
         initial begin
   $display             ("Hello World");



   ;
   ;
       $finish;
end
endmodule
